parameter A_WIDTH = 12;
parameter B_WIDTH = 12;
