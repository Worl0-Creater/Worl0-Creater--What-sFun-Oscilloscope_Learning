`define MODULE_NAME Adder_Subtractor_Top
`define UNSIGNED
`define OVERFLOW
`define ADDER
`define NON_PIPELINE
`define DATA_B
